LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE work.definespack.all;

PACKAGE cupack IS
	CONSTANT base_addr	: positive	:= "4";
	CONSTANT lsb_addr	: positive	:= "5";
	CONSTANT cc_lsb_addr	: positive	:= "6";
	CONSTANT command_len	: positive	:= "23";
	CONSTANT X_IDLE	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0000";
	CONSTANT X_LD_AR	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0001";
	CONSTANT X_LD_AI	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0010";
	CONSTANT X_LD_BR	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0011";
	CONSTANT X_M1	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0100";
	CONSTANT X_M3	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0101";
	CONSTANT X_M2	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0110";
	CONSTANT X_M4	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "0111";
	CONSTANT X_M5	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1000";
	CONSTANT X_M6	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1001";
	CONSTANT X_S5	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1010";
	CONSTANT X_S6	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1011";
	CONSTANT X_RND_BR	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1100";
	CONSTANT X_RND_BI	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1101";
	CONSTANT XS_SND_BI	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1110";
	CONSTANT XC_SND_BI	: std_logic_vector(base_addr-1 DOWNTO 0)	:= "1111";
	CONSTANT S_IDLE	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "100000";
	CONSTANT D_LD_AI	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "000100";
	CONSTANT D_LD_BR	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "000110";
	CONSTANT D_M1	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "001000";
	CONSTANT D_M3	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "001010";
	CONSTANT D_M2	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "001100";
	CONSTANT D_M4	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "001110";
	CONSTANT S_M5	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010000";
	CONSTANT S_M6	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010010";
	CONSTANT S_S5	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010100";
	CONSTANT S_S6	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010110";
	CONSTANT S_RND_BR	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "011000";
	CONSTANT S_RND_BI	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "011010";
	CONSTANT S_SND_BI	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "011100";
	CONSTANT S_LD_AR	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "000011";
	CONSTANT S_LD_AI	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "000101";
	CONSTANT S_LD_BR	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "000111";
	CONSTANT S_M1	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "001001";
	CONSTANT S_M3	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "001011";
	CONSTANT S_M2	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "001101";
	CONSTANT S_M4	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "101111";
	CONSTANT C_M5	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010001";
	CONSTANT C_M6	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010011";
	CONSTANT C_S5	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010101";
	CONSTANT C_S6	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "010111";
	CONSTANT C_RND_BR	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "011001";
	CONSTANT C_RND_BI	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "011011";
	CONSTANT C_SND_BI	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "111101";
	CONSTANT D_IDLE	: std_logic_vector(cc_lsb_addr-1 DOWNTO 0)	:= "100001";
	CONSTANT CW_0	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000000000000000000";
	CONSTANT CW_1	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000100000000000000000";
	CONSTANT CW_2	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00010100000000000000000";
	CONSTANT CW_3	: std_logic_vector(command_len-1 DOWNTO 0)	:= "01001100000000000000000";
	CONSTANT CW_4	: std_logic_vector(command_len-1 DOWNTO 0)	:= "11011101000000000000000";
	CONSTANT CW_5	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00100001000100000000000";
	CONSTANT CW_6	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00100011000110000000000";
	CONSTANT CW_7	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000011100100001100000";
	CONSTANT CW_8	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000001100010001000";
	CONSTANT CW_9	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000010001100001000000";
	CONSTANT CW_10	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000000101110001000";
	CONSTANT CW_11	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000000000001110111";
	CONSTANT CW_12	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000000000000001010";
	CONSTANT CW_13	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000000000000000110";
	CONSTANT CW_14	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000000000000000010";
	CONSTANT CW_15	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000100001100010001000";
	CONSTANT CW_16	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00010110001100001000000";
	CONSTANT CW_17	: std_logic_vector(command_len-1 DOWNTO 0)	:= "01001100000101110001000";
	CONSTANT CW_18	: std_logic_vector(command_len-1 DOWNTO 0)	:= "11011100000000001110111";
	CONSTANT CW_19	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00100000000000000001010";
	CONSTANT CW_20	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00100000000000000000110";
	CONSTANT CW_21	: std_logic_vector(command_len-1 DOWNTO 0)	:= "00000000000000000000010";
END cupack;