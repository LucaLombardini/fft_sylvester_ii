LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE work.definespack.all;

PACKAGE cupack IS
	CONSTANT base_addr	: positive	:= "4";
	CONSTANT lsb_addr	: positive	:= "5";
	CONSTANT cc_lsb_addr	: positive	:= "6";
	CONSTANT command_len	: positive	:= "23";
	CONSTANT uir_width	: positive	:= "29";
	CONSTANT X_IDLE	: std_logic_vector(base_addr-1 DOWNTO 0) := "0000";
	CONSTANT X_LD_AR	: std_logic_vector(base_addr-1 DOWNTO 0) := "0001";
	CONSTANT X_LD_AI	: std_logic_vector(base_addr-1 DOWNTO 0) := "0010";
	CONSTANT X_LD_BR	: std_logic_vector(base_addr-1 DOWNTO 0) := "0011";
	CONSTANT X_M1	: std_logic_vector(base_addr-1 DOWNTO 0) := "0100";
	CONSTANT X_M3	: std_logic_vector(base_addr-1 DOWNTO 0) := "0101";
	CONSTANT X_M2	: std_logic_vector(base_addr-1 DOWNTO 0) := "0110";
	CONSTANT X_M4	: std_logic_vector(base_addr-1 DOWNTO 0) := "0111";
	CONSTANT X_M5	: std_logic_vector(base_addr-1 DOWNTO 0) := "1000";
	CONSTANT X_M6	: std_logic_vector(base_addr-1 DOWNTO 0) := "1001";
	CONSTANT X_S5	: std_logic_vector(base_addr-1 DOWNTO 0) := "1010";
	CONSTANT X_S6	: std_logic_vector(base_addr-1 DOWNTO 0) := "1011";
	CONSTANT X_RND_BR	: std_logic_vector(base_addr-1 DOWNTO 0) := "1100";
	CONSTANT X_RND_BI	: std_logic_vector(base_addr-1 DOWNTO 0) := "1101";
	CONSTANT XS_SND_BI	: std_logic_vector(base_addr-1 DOWNTO 0) := "1110";
	CONSTANT XC_SND_BI	: std_logic_vector(base_addr-1 DOWNTO 0) := "1111";
	CONSTANT IDLE	: std_logic_vector(base_addr-1 DOWNTO 0) := "0000";
	CONSTANT S_LD_AR	: std_logic_vector(base_addr-1 DOWNTO 0) := "0001";
	CONSTANT S_LD_AI	: std_logic_vector(base_addr-1 DOWNTO 0) := "0010";
	CONSTANT S_LD_BR	: std_logic_vector(base_addr-1 DOWNTO 0) := "0011";
	CONSTANT S_M1	: std_logic_vector(base_addr-1 DOWNTO 0) := "0100";
	CONSTANT S_M3	: std_logic_vector(base_addr-1 DOWNTO 0) := "0101";
	CONSTANT S_M2	: std_logic_vector(base_addr-1 DOWNTO 0) := "0110";
	CONSTANT S_M4	: std_logic_vector(base_addr-1 DOWNTO 0) := "0111";
	CONSTANT S_M5	: std_logic_vector(base_addr-1 DOWNTO 0) := "1000";
	CONSTANT S_M6	: std_logic_vector(base_addr-1 DOWNTO 0) := "1001";
	CONSTANT S_S5	: std_logic_vector(base_addr-1 DOWNTO 0) := "1010";
	CONSTANT S_S6	: std_logic_vector(base_addr-1 DOWNTO 0) := "1011";
	CONSTANT S_RND_BR	: std_logic_vector(base_addr-1 DOWNTO 0) := "1100";
	CONSTANT S_RND_BI	: std_logic_vector(base_addr-1 DOWNTO 0) := "1101";
	CONSTANT S_SND_BI	: std_logic_vector(base_addr-1 DOWNTO 0) := "1110";
	CONSTANT C_SND_BI	: std_logic_vector(base_addr-1 DOWNTO 0) := "1111";
	CONSTANT C_M5	: std_logic_vector(base_addr-1 DOWNTO 0) := "1000";
	CONSTANT C_M6	: std_logic_vector(base_addr-1 DOWNTO 0) := "1001";
	CONSTANT C_S5	: std_logic_vector(base_addr-1 DOWNTO 0) := "1010";
	CONSTANT C_S6	: std_logic_vector(base_addr-1 DOWNTO 0) := "1011";
	CONSTANT C_RND_BR	: std_logic_vector(base_addr-1 DOWNTO 0) := "1100";
	CONSTANT C_RND_BI	: std_logic_vector(base_addr-1 DOWNTO 0) := "1101";
	CONSTANT CW_IDLE	: std_logic_vector(command_len-1 DOWNTO 0) := "00000000000000000000000";
	CONSTANT CW_SLD_AR	: std_logic_vector(command_len-1 DOWNTO 0) := "00000100000000000000000";
	CONSTANT CW_SLD_AI	: std_logic_vector(command_len-1 DOWNTO 0) := "00010100000000000000000";
	CONSTANT CW_SLD_BR	: std_logic_vector(command_len-1 DOWNTO 0) := "01001100000000000000000";
	CONSTANT CW_SM1	: std_logic_vector(command_len-1 DOWNTO 0) := "11011101000000000000000";
	CONSTANT CW_SM3	: std_logic_vector(command_len-1 DOWNTO 0) := "00100001000100000000000";
	CONSTANT CW_SM2	: std_logic_vector(command_len-1 DOWNTO 0) := "00100011000110000000000";
	CONSTANT CW_SM4	: std_logic_vector(command_len-1 DOWNTO 0) := "00000011100100001100000";
	CONSTANT CW_SM5	: std_logic_vector(command_len-1 DOWNTO 0) := "00000000001100010001000";
	CONSTANT CW_SM6	: std_logic_vector(command_len-1 DOWNTO 0) := "00000010001100001000000";
	CONSTANT CW_SS5	: std_logic_vector(command_len-1 DOWNTO 0) := "00000000000101110001000";
	CONSTANT CW_SS6	: std_logic_vector(command_len-1 DOWNTO 0) := "00000000000000001110111";
	CONSTANT CW_SRND_BR	: std_logic_vector(command_len-1 DOWNTO 0) := "00000000000000000001010";
	CONSTANT CW_SRND_BI	: std_logic_vector(command_len-1 DOWNTO 0) := "00000000000000000000110";
	CONSTANT CW_SSND_BI	: std_logic_vector(command_len-1 DOWNTO 0) := "00000000000000000000010";
	CONSTANT CW_CM5	: std_logic_vector(command_len-1 DOWNTO 0) := "00000100001100010001000";
	CONSTANT CW_CM6	: std_logic_vector(command_len-1 DOWNTO 0) := "00010110001100001000000";
	CONSTANT CW_CS5	: std_logic_vector(command_len-1 DOWNTO 0) := "01001100000101110001000";
	CONSTANT CW_CS6	: std_logic_vector(command_len-1 DOWNTO 0) := "11011101000000001110111";
	CONSTANT CW_CRND_BR	: std_logic_vector(command_len-1 DOWNTO 0) := "00100001000100000001010";
	CONSTANT CW_CRND_BI	: std_logic_vector(command_len-1 DOWNTO 0) := "00100011000110000000110";
	CONSTANT CW_CSND_BI	: std_logic_vector(command_len-1 DOWNTO 0) := "00000011100100001100010";
END cupack;